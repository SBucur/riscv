import uvm_pkg::*;
`include "uvm_macros.svh"

module test_top();

endmodule