module dut_dummy(
    input clk,
    input rst,
    input [31:0] in_instr,
    input [31:0] in_data,
    output [31:0] pc,
    output [31:0] alu_out,
    output [31:0] out_instr,
    output [31:0] out_data
);

endmodule