`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Author: Stefan Bucur 
// 
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module top(

    );
endmodule
